*INV_Transient_Response
.include TSMC_180nm.txt
.param LAMBDA=0.09u
.param width_P={20*LAMBDA}
.param width_N={10*LAMBDA}
.global gnd vdd


Vdd vdd gnd 1.8V

vin x gnd pulse 0 1.8 0ns 1ns 1ns 10ns 20ns


M1 y x gnd gnd CMOSN W = {width_N} L = {2*LAMBDA}
+ AS = {5*width_N*LAMBDA} PS = {10*LAMBDA + 2*width_N}
+ AD = {5*width_N*LAMBDA} PD = {10*LAMBDA + 2*width_N}

M2 y x vdd vdd CMOSP W = {width_P} L = {2*LAMBDA}
+ AS = {5*width_N*LAMBDA} PS = {10*LAMBDA + 2*width_N}
+ AD = {5*width_N*LAMBDA} PD = {10*LAMBDA + 2*width_N}

Cout y gnd 100f

.tran 0.1n 200n

.control
run 
plot v(y) v(x)
*setting_BG_colour
set color0 = white
set color1 = black
set xbrushwidth = 5
.endc
