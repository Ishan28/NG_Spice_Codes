*MOS_CHAR
.include TSMC_180nm.txt
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.global gnd vdd




VGS G gnd 1.8V
VDS D gnd 1V

M1 D G gnd gnd CMOSN W = {width_N} L = {2*LAMBDA}
+ AS = {5+width_N*LAMBDA} PS = {10*LAMBDA + 2*width_N}
+ AD = {5+width_N*LAMBDA} PD = {10*LAMBDA + 2*width_N}

.dc VGS 0 1.8 0.05

.control
run 
plot -VDS#branch
*setting_BG_colour
set color0 = white
set color1 = black
set xbrushwidth = 5
.endc
